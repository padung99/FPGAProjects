--library ieee;
--use ieee.std_logic_1164.all;
--
--entity test_uart_trans is
--end test_uart_trans;
--
--architecture arch of test_uart_trans is

