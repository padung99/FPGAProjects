library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;


entity instr_mem is
port(
		address: in std_logic_vector(31 downto 0);
		reset: in std_logic;
		o_instr: out std_logic_vector(31 downto 0)
		);
end instr_mem;

architecture arch of instr_mem is

type instruction_memory is array(0 to 31) of std_logic_vector(31 downto 0);
signal RAM: instruction_memory := (
												x"02114020", -------- 0x40 0000 add $t0, $s0, $s1 -- 0000 0010 0001 0001 0100 0000 0010 0000 -- R type
												x"02324822", -------- 0x40 0004 sub $t1, $s1, $s2 -- 0000 0010 0011 0010 0100 1000 0010 0010 -- R type
												x"02115024", -------- 0x40 0008 and $t2, $s0, $s1 -- 0000 0010 0001 0001 0101 0000 0010 0100 -- R type
												x"02535825", -------- 0x40 000C or  $t3, $s2, $s3 -- 0000 0010 0101 0011 0101 1000 0010 0101 -- R type
												x"0211602A", -------- 0x40 0010 slt $t4, $s0, $s1 -- 0000 0010 0001 0001 0110 0000 0010 1010 -- R type
												x"02336820", -------- 0x40 0014 add $t5, $s1, $s3 -- 0000 0010 0011 0011 0110 1000 0010 0000 -- R type
												x"02114020", -------- 0x40 0018 add $t0, $s0, $s1 -- 0000 0010 0001 0001 0100 0000 0010 0000 -- R type
												x"02114020", -------- 0x40 001C add $t0, $s0, $s1 -- 0000 0010 0001 0001 0100 0000 0010 0000 -- R type
												x"02324822", -------- 0x40 0020 sub $t1, $s1, $s2 -- 0000 0010 0011 0010 0100 1000 0010 0010 -- R type
												x"02115024", -------- 0x40 002C slt $t4, $s0, $s1 -- 0000 0010 0001 0001 0110 0000 0010 1010 -- R type
												x"02336820", -------- 0x40 0024 and $t2, $s0, $s1 -- 0000 0010 0001 0001 0101 0000 0010 0100 -- R type
												x"02535825", -------- 0x40 0028 or  $t3, $s2, $s3 -- 0000 0010 0101 0011 0101 1000 0010 0101 -- R type
												x"0211602A", -------- 0x40 0030 add $t5, $s1, $s3 -- 0000 0010 0011 0011 0110 1000 0010 0000 -- R type
												x"02114020", -------- 0x40 0034 add $t0, $s0, $s1 -- 0000 0010 0001 0001 0100 0000 0010 0000 -- R type												
												x"8E280012", -------- 0x40 0038 lw $t0, 12($s1) --   1000 1110 0010 1000 0000 0000 0001 0010 I-type
												x"AE320008", -------- 0x40 003C sw $s2, 8($s1)  --   1010 1110 0011 0010 0000 0000 0000 1000 I_ type
												x"08100008", -------- 0x40 0040 j 0x00400020 -- 0000 1000 0001 0000 0000 0000 0000 1000  -- J type
												
												x"02114020", -------- 0x40 0000 add $t0, $s0, $s1 -- 0000 0010 0001 0001 0100 0000 0010 0000 -- R type
												x"02324822", -------- 0x40 0004 sub $t1, $s1, $s2 -- 0000 0010 0011 0010 0100 1000 0010 0010 -- R type
												x"02115024", -------- 0x40 0008 and $t2, $s0, $s1 -- 0000 0010 0001 0001 0101 0000 0010 0100 -- R type
												x"02535825", -------- 0x40 000C or  $t3, $s2, $s3 -- 0000 0010 0101 0011 0101 1000 0010 0101 -- R type
												x"0211602A", -------- 0x40 0010 slt $t4, $s0, $s1 -- 0000 0010 0001 0001 0110 0000 0010 1010 -- R type
												x"02336820", -------- 0x40 0014 add $t5, $s1, $s3 -- 0000 0010 0011 0011 0110 1000 0010 0000 -- R type
												x"02114020", -------- 0x40 0018 add $t0, $s0, $s1 -- 0000 0010 0001 0001 0100 0000 0010 0000 -- R type
												x"02114020", -------- 0x40 001C add $t0, $s0, $s1 -- 0000 0010 0001 0001 0100 0000 0010 0000 -- R type
												x"02324822", -------- 0x40 0020 sub $t1, $s1, $s2 -- 0000 0010 0011 0010 0100 1000 0010 0010 -- R type
												x"02115024", -------- 0x40 002C slt $t4, $s0, $s1 -- 0000 0010 0001 0001 0110 0000 0010 1010 -- R type
												x"02535825", -------- 0x40 0028 or  $t3, $s2, $s3 -- 0000 0010 0101 0011 0101 1000 0010 0101 -- R type
												x"0211602A", -------- 0x40 0030 add $t5, $s1, $s3 -- 0000 0010 0011 0011 0110 1000 0010 0000 -- R type
												x"02114020", -------- 0x40 0034 add $t0, $s0, $s1 -- 0000 0010 0001 0001 0100 0000 0010 0000 -- R type
												x"08100000", -------- 0x40 0038 j 0x00400000 -- 0000 1000 0001 0000 0000 0000 0000 0000  -- J type
												x"00000000"  -------- 0x40 003C
												);

begin	
	--- address : 0x00400000 = 4194304 
	----  0x003FFFFc = 4194300 -- reset 
o_instr <=  x"00000000" when (reset = '1' or address = x"003FFFFc") else
			   RAM((to_integer(unsigned(address)) - 4194304)/4);
end arch;